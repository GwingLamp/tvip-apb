//------------------------------------------------------------------------------
//  Copyright 2017 Taichi Ishitani
//
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
//
//  http://www.apache.org/licenses/LICENSE-2.0
//
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
//------------------------------------------------------------------------------
`ifndef ${TVIP_NAME}_MACROS_SVH
`define ${TVIP_NAME}_MACROS_SVH

//add parameter below
//`ifndef ${TVIP_NAME}_ADDRESS_WIDTH
//  `define ${TVIP_NAME}_ADDRESS_WIDTH 16
//`endif


`endif
